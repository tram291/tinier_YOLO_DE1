library verilog;
use verilog.vl_types.all;
entity sub_float_tb is
end sub_float_tb;
