library verilog;
use verilog.vl_types.all;
entity tb_multiply is
end tb_multiply;
