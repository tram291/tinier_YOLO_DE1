library verilog;
use verilog.vl_types.all;
entity resize_layer_tb is
end resize_layer_tb;
