library verilog;
use verilog.vl_types.all;
entity float_convert_tb is
end float_convert_tb;
