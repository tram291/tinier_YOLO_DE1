library verilog;
use verilog.vl_types.all;
entity upsample_controller_tb is
end upsample_controller_tb;
