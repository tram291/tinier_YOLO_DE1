library verilog;
use verilog.vl_types.all;
entity add_float_tb is
end add_float_tb;
