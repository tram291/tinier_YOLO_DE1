library verilog;
use verilog.vl_types.all;
entity reorg_layer_tb is
end reorg_layer_tb;
