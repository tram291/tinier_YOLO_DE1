library verilog;
use verilog.vl_types.all;
entity tb_float_larger is
end tb_float_larger;
