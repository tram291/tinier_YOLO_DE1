module get_box_coord ();
  
endmodule