library verilog;
use verilog.vl_types.all;
entity decimal_extract_tb is
end decimal_extract_tb;
