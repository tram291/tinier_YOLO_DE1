//this module will resize 640x480 to 384x384
`include "parameters.h"
module resize_controller(
    clk,
    reset_n,
    enable,
    src_addr1, 
    src_addr2,
    des_addr,
    stage_flag, 
    fraction_part,
    done
);

  parameter SRC_WIDTH       = 640;
  parameter SRC_HEIGHT      = 480;
  parameter SRC_DEPTH       = 3;
  parameter DES_WIDTH       = 384;
  parameter DES_HEIGHT      = 384;
  parameter WIDTH_SCALE     = 16'h3EAC;  //(640-1)/(384-1)=1.6684 
  parameter HEIGHT_SCALE    = 16'h3D00;  //(480-1)/(384-1)=1.2506

  input wire clk;
  input wire reset_n;
  input wire enable;
  

  output reg  done, stage_flag;
  output reg  [`ADDR_SZ-1:0] src_addr1, src_addr2;
  output reg  [`ADDR_SZ-1:0] des_addr; 
  output wire [15:0] fraction_part;
  
  reg [15:0] row, column;
  reg [15:0] channel;
    
  wire [15:0] w_int_val, w_index, fw_index, fw_int_val, fw_scale; 
  wire [15:0] fw_product;
      
  assign w_index  = stage_flag ? row : column;
  assign fw_scale = stage_flag ? HEIGHT_SCALE : WIDTH_SCALE;
  
  float_convert fc1 (.d(w_index), .f(fw_index));
  Multiply      m1  (.a(fw_scale), .b(fw_index), .result(fw_product)); 
  
  decimal_extract de  (.in(fw_product), .out(w_int_val));  
  float_convert   fc2 (.d(w_int_val), .f(fw_int_val));
  sub_float       sf  (.a(fw_product), .b(fw_int_val), .c(fraction_part));
    

  always @(posedge clk or negedge reset_n) begin
      if (~reset_n) begin
          row           <= 0;
          column        <= 0;
          channel       <= 0;
          src_addr1     <= 0;
          src_addr2     <= 0;
          des_addr      <= 0;
          done          <= 0;
          stage_flag    <= 0;
      end
      else begin
          if (enable & ~done) begin
              if (~stage_flag) begin 
                  column = column + 1;   
                  if (column == DES_WIDTH) begin
                      column = 0;
                      row = row + 1;
                  end
                  if (row == SRC_HEIGHT) begin 
                      row = 0;
                      channel = channel + 1;
                  end 
                  if (channel == SRC_DEPTH) begin
                      channel = 0;
                      stage_flag = 1;
                  end
                  
                  src_addr1 = w_int_val + SRC_WIDTH*(row + SRC_HEIGHT*channel);
                  src_addr2 = src_addr1 + 1;
                  
                  des_addr = column + DES_WIDTH*(row + SRC_HEIGHT*channel);
              end
              else begin                            
                  column = column + 1;
                  if (column > DES_WIDTH) begin
                      column = 0;
                      row = row + 1;
                  end
                  if (row == DES_HEIGHT) begin 
                      row = 0;
                      channel = channel + 1;
                  end 
                  if (channel == SRC_DEPTH) begin
                      channel = 0;
                      done = 1;
                  end
                  
                  src_addr1 = column + DES_WIDTH*(w_int_val + SRC_HEIGHT*channel);
                  src_addr2 = src_addr1 + DES_WIDTH;
                  
                  des_addr = column + DES_WIDTH*(row + DES_HEIGHT*channel);
              end
          end
      end
  end


  
endmodule
