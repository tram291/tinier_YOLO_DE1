library verilog;
use verilog.vl_types.all;
entity tb_resize_datapath is
end tb_resize_datapath;
