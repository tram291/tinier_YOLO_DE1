library verilog;
use verilog.vl_types.all;
entity resize_controller_tb is
end resize_controller_tb;
